library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

entity Timer is
	port (Clock, Start : in std_logic;
		    Data_in : in std_logic_vector(9 downto 0);
		    Time_out : out std_logic;
		    -- Comment out the next 2 lines for running on board.
		    OSeg0, OSeg1, OSeg2 : out std_logic_vector(7 downto 0);
		    OTens_seconds : out std_logic_vector(3 downto 0));
end entity Timer;

architecture arc of Timer is
	component BCD_Counter is
		port (Clk, Direction, Init, Enable : in std_logic;
				  Q_Out : out std_logic_vector(3 downto 0));
	end component BCD_Counter;
	
	component BCD_Counter_Min is
		port (Clk, Direction, Init, Enable : in std_logic;
				  Q_Out : out std_logic_vector(3 downto 0));
	end component BCD_Counter_Min;
	
signal Direction, Init : std_logic;
signal Ones_seconds, Tens_seconds, Minutes : std_logic_vector(3 downto 0);
signal Clock2, Clock3 : std_logic;
signal Seg0, Seg1, Seg2 : std_logic_vector(7 downto 0);
		
begin
  BCD1: BCD_Counter 
    port map (Clk => Clock, Direction => Direction, Init => Init, Enable => Start, Q_Out => Ones_seconds);
      
  BCD2: BCD_Counter_Min
    port map (Clk => Clock2, Direction => Direction, Init => Init, Enable => Start, Q_Out => Tens_seconds);
      
  BCD3: BCD_Counter
    port map (Clk => Clock3, Direction => Direction, Init => Init, Enable => Start, Q_Out => Minutes);
      
  Clock2 <= '1' when Ones_seconds = "0000"
                else '0';
                  
  Clock3 <= '1' when Tens_seconds = "0000"
                else '0';
  
	Direction <= '0';
	Init <= '1';
	
    process (Clock)
    begin
        if RISING_EDGE(Clock) then
           if (Start = '1') then
             
             if ((Minutes = Data_in(9 downto 8)) and (Tens_seconds = Data_in(7 downto 4)) and (Ones_seconds = Data_in(3 downto 0))) then
               Time_out <= '1';
             end if;
             
                case Minutes is
                    when "0000" => Seg0 <= "00000011"; --0
                    when "0001" => Seg0 <= "10011111"; --1
                    when "0010" => Seg0 <= "00100101"; --2
                    when "0011" => Seg0 <= "00001101"; --3
                    when others => Seg0 <= "11111111";
                end case;
                
                case Tens_seconds is
                    when "0000" => Seg1 <= "00000011"; --0
                    when "0001" => Seg1 <= "10011111"; --1
                    when "0010" => Seg1 <= "00100101"; --2
                    when "0011" => Seg1 <= "00001101"; --3
                    when "0100" => Seg1 <= "10011001"; --4
                    when "0101" => Seg1 <= "01001001"; --5
                    when others => Seg1 <= "11111111";
                end case;
                
                case Ones_seconds is
                    when "0000" => Seg2 <= "00000011"; --0
                    when "0001" => Seg2 <= "10011111"; --1
                    when "0010" => Seg2 <= "00100101"; --2
                    when "0011" => Seg2 <= "00001101"; --3
                    when "0100" => Seg2 <= "10011001"; --4
                    when "0101" => Seg2 <= "01001001"; --5
                    when "0110" => Seg2 <= "01000001"; --6
                    when "0111" => Seg2 <= "00011111"; --7
                    when "1000" => Seg2 <= "00000001"; --8
                    when "1001" => Seg2 <= "00001001"; --9
                    when others => Seg2 <= "11111111";
                end case;
                
            else
                Seg0 <= "11111111";
                Seg1 <= "11111111";
                Seg2 <= "11111111";
            end if;
        end if;
    end process;
    
    -- Comment out these lines for running on board.
    OSeg0 <= Seg0;
    OSeg1 <= Seg1;
    OSeg2 <= Seg2;
    OTens_seconds <= Tens_seconds;

end architecture arc;