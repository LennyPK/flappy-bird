library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity ROM is
    port (  address : in integer;
            data    : out integer;
         );
end entity ROM;

architecture behaviour of ROM is
    type mem is array (0 to 99) of integer;
    constant my_rom : mem := (
        -- binary
        -- 00 => "00000000";
        -- 01 => "00000001";
        -- 02 => "00000010";
        -- 03 => "00000011";
        -- 04 => "00000100";
        -- 05 => "00000101";
        -- 06 => "00000110";
        -- 07 => "00000111";
        -- 08 => "00001000";
        -- 09 => "00001001";
        -- 10 => "00001010";
        -- 11 => "00001011";
        -- 12 => "00001100";
        -- 13 => "00001101";
        -- 14 => "00001110";
        -- 15 => "00001111";
        -- 16 => "00010000";
        -- 17 => "00010001";
        -- 18 => "00010010";
        -- 19 => "00010011";
        -- 20 => "00010100";
        -- 21 => "00010101";
        -- 22 => "00010110";
        -- 23 => "00010111";
        -- 24 => "00011000";
        -- 25 => "00011001";
        -- 26 => "00011010";
        -- 27 => "00011011";
        -- 28 => "00011100";
        -- 29 => "00011101";
        -- 30 => "00011110";
        -- 31 => "00011111";
        -- 32 => "00100000";
        -- 33 => "00100001";
        -- 34 => "00100010";
        -- 35 => "00100011";
        -- 36 => "00100100";
        -- 37 => "00100101";
        -- 38 => "00100110";
        -- 39 => "00100111";
        -- 40 => "00101000";
        -- 40 => "00101000";
        -- 41 => "00101001";
        -- 42 => "00101010";
        -- 43 => "00101011";
        -- 44 => "00101100";
        -- 45 => "00101101";
        -- 46 => "00101110";
        -- 47 => "00101111";
        -- 48 => "00110000";
        -- 49 => "00110001";
        -- 50 => "00110010";
        -- 51 => "00110011";
        -- 52 => "00110100";
        -- 53 => "00110101";
        -- 54 => "00110110";
        -- 55 => "00110111";
        -- 56 => "00111000";
        -- 57 => "00111001";
        -- 58 => "00111010";
        -- 59 => "00111011";
        -- 60 => "00111100";
        -- 61 => "00111101";
        -- 62 => "00111110";
        -- 63 => "00111111";
        -- 64 => "01000000";
        -- 65 => "01000001";
        -- 66 => "01000010";
        -- 67 => "01000011";
        -- 68 => "01000100";
        -- 69 => "01000101";
        -- 70 => "01000110";
        -- 71 => "01000111";
        -- 72 => "01001000";
        -- 73 => "01001001";
        -- 74 => "01001010";
        -- 75 => "01001011";
        -- 76 => "01001100";
        -- 77 => "01001101";
        -- 78 => "01001110";
        -- 79 => "01001111";
        -- 80 => "01010000";
        -- 81 => "01010001";
        -- 82 => "01010010";
        -- 83 => "01010011";
        -- 84 => "01010100";
        -- 85 => "01010101";
        -- 86 => "01010110";
        -- 87 => "01010111";
        -- 88 => "01011000";
        -- 89 => "01011001";
        -- 90 => "01011010";
        -- 91 => "01011011";
        -- 92 => "01011100";
        -- 93 => "01011101";
        -- 94 => "01011110";
        -- 95 => "01011111";
        -- 96 => "01100000";
        -- 97 => "01100001";
        -- 98 => "01100010";
        -- 99 => "01100011";

        -- integers
        00 => 00;
        01 => 01;
        02 => 02;
        03 => 03;
        04 => 04;
        05 => 05;
        06 => 06;
        07 => 07;
        08 => 08;
        09 => 09;
        10 => 10;
        11 => 11;
        12 => 12;
        13 => 13;
        14 => 14;
        15 => 15;
        16 => 16;
        17 => 17;
        18 => 18;
        19 => 19;
        20 => 20;
        21 => 21;
        22 => 22;
        23 => 23;
        24 => 24;
        25 => 25;
        26 => 26;
        27 => 27;
        28 => 28;
        29 => 29;
        30 => 30;
        31 => 31;
        32 => 32;
        33 => 33;
        34 => 34;
        35 => 35;
        36 => 36;
        37 => 37;
        38 => 38;
        39 => 39;
        40 => 40;
        41 => 41;
        42 => 42;
        43 => 43;
        44 => 44;
        45 => 45;
        46 => 46;
        47 => 47;
        48 => 48;
        49 => 49;
        50 => 50;
        51 => 51;
        52 => 52;
        53 => 53;
        54 => 54;
        55 => 55;
        56 => 56;
        57 => 57;
        58 => 58;
        59 => 59;
        60 => 60;
        61 => 61;
        62 => 62;
        63 => 63;
        64 => 64;
        65 => 65;
        66 => 66;
        67 => 67;
        68 => 68;
        69 => 69;
        70 => 70;
        71 => 71;
        72 => 72;
        73 => 73;
        74 => 74;
        75 => 75;
        76 => 76;
        77 => 77;
        78 => 78;
        79 => 79;
        80 => 80;
        81 => 81;
        82 => 82;
        83 => 83;
        84 => 84;
        85 => 85;
        86 => 86;
        87 => 87;
        88 => 88;
        89 => 89;
        90 => 90;
        91 => 91;
        92 => 92;
        93 => 93;
        94 => 94;
        95 => 95;
        96 => 96;
        97 => 97;
        98 => 98;
        99 => 99;
    );
begin
    process (address)
    begin
        case address is
            when 0 => data <= my_rom(0);
            when 1 => data <= my_rom(1);
            when 2 => data <= my_rom(2);
            when 3 => data <= my_rom(3);
            when 4 => data <= my_rom(4);
            when 5 => data <= my_rom(5);
            when 6 => data <= my_rom(6);
            when 7 => data <= my_rom(7);
            when 8 => data <= my_rom(8);
            when 9 => data <= my_rom(9);
            when 10 => data <= my_rom(10);
            when 11 => data <= my_rom(11);
            when 12 => data <= my_rom(12);
            when 13 => data <= my_rom(13);
            when 14 => data <= my_rom(14);
            when 15 => data <= my_rom(15);
            when 16 => data <= my_rom(16);
            when 17 => data <= my_rom(17);
            when 18 => data <= my_rom(18);
            when 19 => data <= my_rom(19);
            when 20 => data <= my_rom(20);
            when 21 => data <= my_rom(21);
            when 22 => data <= my_rom(22);
            when 23 => data <= my_rom(23);
            when 24 => data <= my_rom(24);
            when 25 => data <= my_rom(25);
            when 26 => data <= my_rom(26);
            when 27 => data <= my_rom(27);
            when 28 => data <= my_rom(28);
            when 29 => data <= my_rom(29);
            when 30 => data <= my_rom(30);
            when 31 => data <= my_rom(31);
            when 32 => data <= my_rom(32);
            when 33 => data <= my_rom(33);
            when 34 => data <= my_rom(34);
            when 35 => data <= my_rom(35);
            when 36 => data <= my_rom(36);
            when 37 => data <= my_rom(37);
            when 38 => data <= my_rom(38);
            when 39 => data <= my_rom(39);
            when 40 => data <= my_rom(40);
            when 41 => data <= my_rom(41);
            when 42 => data <= my_rom(42);
            when 43 => data <= my_rom(43);
            when 44 => data <= my_rom(44);
            when 45 => data <= my_rom(45);
            when 46 => data <= my_rom(46);
            when 47 => data <= my_rom(47);
            when 48 => data <= my_rom(48);
            when 49 => data <= my_rom(49);
            when 50 => data <= my_rom(50);
            when 51 => data <= my_rom(51);
            when 52 => data <= my_rom(52);
            when 53 => data <= my_rom(53);
            when 54 => data <= my_rom(54);
            when 55 => data <= my_rom(55);
            when 56 => data <= my_rom(56);
            when 57 => data <= my_rom(57);
            when 58 => data <= my_rom(58);
            when 59 => data <= my_rom(59);
            when 60 => data <= my_rom(60);
            when 61 => data <= my_rom(61);
            when 62 => data <= my_rom(62);
            when 63 => data <= my_rom(63);
            when 64 => data <= my_rom(64);
            when 65 => data <= my_rom(65);
            when 66 => data <= my_rom(66);
            when 67 => data <= my_rom(67);
            when 68 => data <= my_rom(68);
            when 69 => data <= my_rom(69);
            when 70 => data <= my_rom(70);
            when 71 => data <= my_rom(71);
            when 72 => data <= my_rom(72);
            when 73 => data <= my_rom(73);
            when 74 => data <= my_rom(74);
            when 75 => data <= my_rom(75);
            when 76 => data <= my_rom(76);
            when 77 => data <= my_rom(77);
            when 78 => data <= my_rom(78);
            when 79 => data <= my_rom(79);
            when 80 => data <= my_rom(80);
            when 81 => data <= my_rom(81);
            when 82 => data <= my_rom(82);
            when 83 => data <= my_rom(83);
            when 84 => data <= my_rom(84);
            when 85 => data <= my_rom(85);
            when 86 => data <= my_rom(86);
            when 87 => data <= my_rom(87);
            when 88 => data <= my_rom(88);
            when 89 => data <= my_rom(89);
            when 90 => data <= my_rom(90);
            when 91 => data <= my_rom(91);
            when 92 => data <= my_rom(92);
            when 93 => data <= my_rom(93);
            when 94 => data <= my_rom(94);
            when 95 => data <= my_rom(95);
            when 96 => data <= my_rom(96);
            when 97 => data <= my_rom(97);
            when 98 => data <= my_rom(98);
            when 99 => data <= my_rom(99);
        end case;
    end process;
end architecture behaviour;
